library verilog;
use verilog.vl_types.all;
entity isgreater_64bit_vlg_vec_tst is
end isgreater_64bit_vlg_vec_tst;
