library verilog;
use verilog.vl_types.all;
entity DATAPATH_vlg_vec_tst is
end DATAPATH_vlg_vec_tst;
