library verilog;
use verilog.vl_types.all;
entity and_self_vlg_vec_tst is
end and_self_vlg_vec_tst;
