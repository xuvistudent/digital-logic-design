module full_sub_32bit(	input [31:0] a,
								input [31:0] b,
								input c_in,
								output c_out,
								output [31:0] res);
	assign {c_out, res} = a + ~b + c_in;
endmodule