module and_1bit(	input a,
						input b,
						output c);
	assign c = a & b;
endmodule