library verilog;
use verilog.vl_types.all;
entity set_bit_0_vlg_vec_tst is
end set_bit_0_vlg_vec_tst;
